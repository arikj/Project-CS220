module FA(input a,b, cin, output wire sum );

xor x1(sum, a, b, cin);

endmodule
